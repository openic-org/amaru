** sch_path: /home/designer/shared/amaru/analog/tb/tb_lskmod_gen.sch
**.subckt tb_lskmod_gen
V2 VSS GND 0
V1 VG VSS 0
I0 VIP VIN dc 0 ac 1
C2 VIP VIN 2.72p m=1
L1 net1 VIN 47n m=1
R1 VIP net1 0.471 m=1
C1 VIP VIN 0.15412p m=1
XM2 VIN VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM3 VIP VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
x1 VIP VSS VG VIN lskmod_py_47e-9_0_471_1870e6_289_433e6
**** begin user architecture code


.lib cornerMOSlv.lib mos_tt





.save all
.save V(VIP) V(VIN)
.ac dec 1000 350Meg 550Meg

.control
  set filetype=ascii        ; ASCII .raw (human-readable)
  run
  alter v1 dc=1.2
  run
  let ZIN0  = ac1.v(VIP) - ac1.v(VIN)
  let ABSZ0 = abs(ZIN0)
  let IMZ0  = imag(ZIN0)
  let REZ0  = real(ZIN0)
  let Q0    = IMZ0/REZ0
  let ZIN1  = ac2.v(VIP) - ac2.v(VIN)
  let ABSZ1 = abs(ZIN1)
  let IMZ1  = imag(ZIN1)
  let REZ1  = real(ZIN1)
  let Q1    = IMZ1/REZ1
  write tb_lskm_g1.raw ABSZ0 Q0 ABSZ1 Q1
  set appendwrite
.endc


**** end user architecture code
**.ends

* expanding   symbol:  lskmod_gen.sym # of pins=4
** sym_path: /home/designer/shared/amaru/analog/core/lskmod_gen.sym
** sch_path: /home/designer/shared/amaru/analog/core/lskmod_gen.sch
.subckt lskmod_gen VA VSS D VB
*.iopin VA
*.iopin VSS
*.iopin D
*.iopin VB
XM1 VA D VB VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  lskmod.py(47e-9,0.471,1870e6,289,433e6) # of pins=4
** sym_path: /home/designer/shared/amaru/analog/core/lskmod_gen.sym
** sch_path: /home/designer/shared/amaru/analog/core/lskmod.py
.subckt lskmod_py_47e-9_0_471_1870e6_289_433e6 VA VSS D VB
*.iopin VA
*.iopin VSS
*.iopin D
*.iopin VB
XM1 VA D VB VSS sg13_lv_nmos w=3.91u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
