** sch_path: /home/designer/shared/amaru/analog/tb/tb_coil.sch
**.subckt tb_coil
L1 net1 VIN 100n m=1
R1 VIP net1 0.34 m=1
C1 VIP VIN 0.39578p m=1
V17 VSS GND 0
R2 VIP VSS 75k m=1
R3 VSS VIN 75k m=1
I0 VIP VIN dc 0 ac 1
**** begin user architecture code



.save all
.save V(VIP) V(VIN) V(VIP, VIN)
.save I(VPORT)


.control
  set filetype=ascii        ; ASCII .raw (human-readable)
    run
    ac dec 1000 1Meg 1000Meg
    *tran 0.1u 100u
    let ZIN  = v(VIP, VIN)
    let ABSZ = abs(ZIN)
    let IMZ  = imag(ZIN)
    let REZ  = real(ZIN)
    let Q    = IMZ/REZ
    meas ac F_res when IMZ=0
    write tb_coil1.raw ABSZ Q
    set appendwrite
.endc



.lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
