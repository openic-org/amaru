** sch_path: /home/designer/shared/amaru/analog/tb/tb_ldo_01_stb.sch
**.subckt tb_ldo_01_stb
C1 VLDO VSS 253.58n m=1
V1 VDD GND 1.3
V2 VSS GND 0
V3 VREF VSS 0.6
x1 VDD net1 net3 VSS VREF opamp_01
XM1 VLDO net3 VDD VDD sg13_lv_pmos w=91.33u l=0.5u ng=10 m=1
R2 net2 VSS 500k m=1
R1 VLDO net2 500k m=1
R3 VLDO VSS 240k m=1
X999 net1 net2 loopgainprobe
**** begin user architecture code


.param temp=27
.options savecurrents
.ac dec 80 1 10g
.save all v(X999.x) i(v.X999.Vi)
+ @n.xm1.nsg13_lv_pmos[ids]
+ @n.xm1.nsg13_lv_pmos[gm]
+ @n.xm1.nsg13_lv_pmos[gds]

.control
  run
  alter i.X999.Ii acmag=1
  alter v.X999.Vi acmag=0
  run

  let A=ac2.i(v.X999.Vi)
  let B=ac1.i(v.X999.Vi)
  let C=ac2.v(X999.x)
  let D=ac1.v(X999.x)
  let Ttian=(2*(B*C-A*D)+D+A)/(2*(B*C-A*D)+A+D-1)

  set filetype=ascii
  write tb_ldo_02_stb.raw db(Ttian) 180*cph(Ttian)/pi

  set appendwrite
  op
  set filetype=ascii
  write tb_ldo_01_op_stb.raw
.endc




.lib cornerMOSlv.lib mos_tt


**** end user architecture code
**.ends

* expanding   symbol:  opamp_01.sym # of pins=5
** sym_path: /home/designer/shared/amaru/analog/core/opamp_01.sym
** sch_path: /home/designer/shared/amaru/analog/core/opamp_01.sch
.subckt opamp_01 VDD VIP VO VSS VIM
*.iopin VIM
*.iopin VIP
*.iopin VSS
*.iopin VDD
*.iopin VO
XM1 net2 VIP net1 VSS sg13_lv_nmos w=10u l=0.25u ng=1 m=1
XM2 VO VIM net1 VSS sg13_lv_nmos w=10u l=0.25u ng=1 m=1
XM3 net2 net2 VDD VDD sg13_lv_pmos w=1u l=4u ng=1 m=1
XM4 VO net2 VDD VDD sg13_lv_pmos w=1u l=4u ng=1 m=1
XM5 net1 net3 VSS VSS sg13_lv_nmos w=2u l=2u ng=1 m=1
XM6 net3 net3 VSS VSS sg13_lv_nmos w=2u l=2u ng=1 m=1
I0 VDD net3 100n
.ends


* expanding   symbol:  loopgainprobe.sym # of pins=2
** sym_path: /home/designer/shared/amaru/analog/tb/loopgainprobe.sym
** sch_path: /home/designer/shared/amaru/analog/tb/loopgainprobe.sch
.subckt loopgainprobe b a
*.iopin a
*.iopin b
Vi x a dc 0 ac 1
Ii GND x dc 0 ac 0
Vnodebuffer b x 0
.ends

.GLOBAL GND
.end
