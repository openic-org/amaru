* Extracted by KLayout with SG13G2 LVS runset on : 23/08/2025 11:42

.SUBCKT inv_1x VSS Z A VDD
M$1 VSS A Z VSS sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$2 VDD A Z VDD sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u PD=4.68u
.ENDS inv_1x
