** sch_path: /home/designer/shared/amaru/analog/tb/tb_ldo_01.sch
**.subckt tb_ldo_01
C1 VLDO VSS 253.58n m=1
V1 VDD GND dc 1.3 ac 1
V2 VSS GND 0
V3 VREF VSS 0.6
x1 VDD net1 net2 VSS VREF opamp_01
XM1 VLDO net2 VDD VDD sg13_lv_pmos w=91.33u l=0.5u ng=10 m=1
R2 net1 VSS 500k m=1
R1 VLDO net1 500k m=1
R3 VLDO VSS 240k m=1
**** begin user architecture code


.param temp=27
.options savecurrents
.op
.save all
+ @n.xm1.nsg13_lv_pmos[ids]
+ @n.xm1.nsg13_lv_pmos[gm]
+ @n.xm1.nsg13_lv_pmos[gds]

.control
  ac dec 160 10 1g
  set filetype=ascii
  set units=degress
  let PSRR = 1/VLDO
  write tb_ldo_02.raw vdb(PSRR) vp(PSRR)
  set appendwrite
.endc




.lib cornerMOSlv.lib mos_tt


**** end user architecture code
**.ends

* expanding   symbol:  opamp_01.sym # of pins=5
** sym_path: /home/designer/shared/amaru/analog/core/opamp_01.sym
** sch_path: /home/designer/shared/amaru/analog/core/opamp_01.sch
.subckt opamp_01 VDD VIP VO VSS VIM
*.iopin VIM
*.iopin VIP
*.iopin VSS
*.iopin VDD
*.iopin VO
XM1 net2 VIP net1 VSS sg13_lv_nmos w=10u l=0.25u ng=1 m=1
XM2 VO VIM net1 VSS sg13_lv_nmos w=10u l=0.25u ng=1 m=1
XM3 net2 net2 VDD VDD sg13_lv_pmos w=1u l=4u ng=1 m=1
XM4 VO net2 VDD VDD sg13_lv_pmos w=1u l=4u ng=1 m=1
XM5 net1 net3 VSS VSS sg13_lv_nmos w=2u l=2u ng=1 m=1
XM6 net3 net3 VSS VSS sg13_lv_nmos w=2u l=2u ng=1 m=1
I0 VDD net3 100n
.ends

.GLOBAL GND
.end
