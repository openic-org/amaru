** sch_path: /home/designer/shared/amaru/analog/tb/tb_nmos_lv_vgs.sch
**.subckt tb_nmos_lv_vgs
V1 VDD GND 0.75
V2 VSS GND 0
V3 VG GND 0.75
XM1 VDD VG VSS VSS sg13_lv_nmos w=widthn l=lengthn ng=1 m=1
**** begin user architecture code


.param temp=27
.param widthn=1u
.param lengthn=0.5u
.dc v3 0 1.5 0.01
.save @n.xm1.nsg13_lv_nmos[ids]
.save @n.xm1.nsg13_lv_nmos[vth]
.save @n.xm1.nsg13_lv_nmos[gm]
.save @n.xm1.nsg13_lv_nmos[gmb]
.save @n.xm1.nsg13_lv_nmos[gds]
.save @n.xm1.nsg13_lv_nmos[cgg]
.save @n.xm1.nsg13_lv_nmos[cgs]
.save @n.xm1.nsg13_lv_nmos[cgd]
.save @n.xm1.nsg13_lv_nmos[cgb]
.save @n.xm1.nsg13_lv_nmos[cdd]
.save @n.xm1.nsg13_lv_nmos[css]
.save @n.xm1.nsg13_lv_nmos[cgsol]
.save @n.xm1.nsg13_lv_nmos[cgdol]
.save @n.xm1.nsg13_lv_nmos[cjs]
.save @n.xm1.nsg13_lv_nmos[cjd]

.control
  set filetype = ascii
  foreach wval 10u 50u 200u 500u
    alterparam widthn = $wval
    reset
    run
    let ids = @n.xm1.nsg13_lv_nmos[ids]
    let vth = @n.xm1.nsg13_lv_nmos[vth]
    let gm = @n.xm1.nsg13_lv_nmos[gm]
    let gmb = @n.xm1.nsg13_lv_nmos[gmb]
    let gds = @n.xm1.nsg13_lv_nmos[gds]
    let cgg = @n.xm1.nsg13_lv_nmos[cgg]
    let cgs = @n.xm1.nsg13_lv_nmos[cgs]
    let cgd = @n.xm1.nsg13_lv_nmos[cgd]
    let cgb = @n.xm1.nsg13_lv_nmos[cgb]
    let cdd = @n.xm1.nsg13_lv_nmos[cdd]
    let css = @n.xm1.nsg13_lv_nmos[css]
    let cgsol = @n.xm1.nsg13_lv_nmos[cgsol]
    let cgdol = @n.xm1.nsg13_lv_nmos[cgdol]
    let cjs = @n.xm1.nsg13_lv_nmos[cjs]
    let cjd = @n.xm1.nsg13_lv_nmos[cjd]
    write nmoslv_vgs2.raw ids vth gm gmb gds cgg cgs cgd cgb cdd css cgsol cgdol cjs cjd
    set appendwrite
  end
.endc





.lib cornerMOSlv.lib mos_tt


**** end user architecture code
**.ends
.GLOBAL GND
.end
