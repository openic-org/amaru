** sch_path: /home/designer/shared/amaru/analog/tb/tb_nmos_lv_vds.sch
**.subckt tb_nmos_lv_vds
V1 VDD GND 0.75
V2 VSS GND 0
V3 VG GND 0.75
XM1 VDD VG VSS VSS sg13_lv_nmos w=widthn l=lengthn ng=1 m=1
**** begin user architecture code


.param temp=27
.param widthn=1u
.param lengthn=1u
.dc v1 0 1.5 0.01
.save @n.xm1.nsg13_lv_nmos[ids]

.control
  set filetype = ascii
  foreach wval 10u 50u 200u 500u
    alterparam widthn = $wval
    reset
    run
    let ids = @n.xm1.nsg13_lv_nmos[ids]
    let ro = 1/deriv(ids)
    write nmoslv_vds3.raw ids ro
    set appendwrite
  end
.endc





.lib cornerMOSlv.lib mos_tt


**** end user architecture code
**.ends
.GLOBAL GND
.end
