** sch_path: /home/designer/shared/amaru/analog/tb/tb_ldo_gen_stb_2.sch
**.subckt tb_ldo_gen_stb_2
V1 VDD GND 1.2
V2 VSS GND 0
V3 VREF VSS 0.6
R3 VLDO VSS 183.33k m=1
X999 net2 net1 loopgainprobe
x1 VREF VLDO net2 VSS net1 VDD ldo01_py_6e-6_1_1_1_2_0_6
**** begin user architecture code


.param temp=27
.options savecurrents
.ac dec 80 1 10g
.save all v(X999.x) i(v.X999.Vi)
+ @n.x1.xm1.nsg13_lv_pmos[ids]
+ @n.x1.xm1.nsg13_lv_pmos[gm]
+ @n.x1.xm1.nsg13_lv_pmos[gds]

.control
  run
  alter i.X999.Ii acmag=1
  alter v.X999.Vi acmag=0
  run

  let A=ac2.i(v.X999.Vi)
  let B=ac1.i(v.X999.Vi)
  let C=ac2.v(X999.x)
  let D=ac1.v(X999.x)
  let Ttian=(2*(B*C-A*D)+D+A)/(2*(B*C-A*D)+A+D-1)

  set filetype=ascii
  write tb_ldo_g2_stb.raw db(Ttian) 180*cph(Ttian)/pi

  set appendwrite
  op
  set filetype=ascii
  write tb_ldo_gen_stb2.raw
.endc




.lib cornerMOSlv.lib mos_tt


**** end user architecture code
**.ends

* expanding   symbol:  loopgainprobe.sym # of pins=2
** sym_path: /home/designer/shared/amaru/analog/tb/loopgainprobe.sym
** sch_path: /home/designer/shared/amaru/analog/tb/loopgainprobe.sch
.subckt loopgainprobe b a
*.iopin a
*.iopin b
Vi x a dc 0 ac 1
Ii GND x dc 0 ac 0
Vnodebuffer b x 0
.ends


* expanding   symbol:  ldo_01_gen.sym # of pins=6
** sym_path: /home/designer/shared/amaru/analog/core/ldo_01_gen.sym
** sch_path: /home/designer/shared/amaru/analog/core/ldo_01_gen.sch
.subckt ldo_01_gen VREF VLDO VB VSS VA VDD
*.iopin VREF
*.iopin VLDO
*.iopin VDD
*.iopin VB
*.iopin VSS
*.iopin VA
C1 VLDO VSS 1n m=1
x1 VDD VB VG VSS VREF opamp_01
XM1 VLDO VG VDD VDD sg13_lv_pmos w=1u l=0.13u ng=1 m=1
R2 VA VSS 500k m=1
R1 VLDO VA 500k m=1
.ends


* expanding   symbol:  ldo01.py(6e-6,1.1,1.2,0.6) # of pins=6
** sym_path: /home/designer/shared/amaru/analog/core/ldo_01_gen.sym
** sch_path: /home/designer/shared/amaru/analog/core/ldo01.py
.subckt ldo01_py_6e-6_1_1_1_2_0_6 VREF VLDO VB VSS VA VDD
*.iopin VREF
*.iopin VLDO
*.iopin VDD
*.iopin VB
*.iopin VSS
*.iopin VA
C1 VLDO VSS 19.16n m=1
R1 VLDO VA 416.67k m=1
R2 VA VSS 500.0k m=1
XM1 VLDO VG VDD VDD sg13_lv_pmos w=14.84u l=0.25u ng=2 m=1
x1 VDD VB VG VSS VREF opamp_01
.ends


* expanding   symbol:  opamp_01.sym # of pins=5
** sym_path: /home/designer/shared/amaru/analog/core/opamp_01.sym
** sch_path: /home/designer/shared/amaru/analog/core/opamp_01.sch
.subckt opamp_01 VDD VIP VO VSS VIM
*.iopin VIM
*.iopin VIP
*.iopin VSS
*.iopin VDD
*.iopin VO
XM1 net2 VIP net1 VSS sg13_lv_nmos w=10u l=0.25u ng=1 m=1
XM2 VO VIM net1 VSS sg13_lv_nmos w=10u l=0.25u ng=1 m=1
XM3 net2 net2 VDD VDD sg13_lv_pmos w=1u l=4u ng=1 m=1
XM4 VO net2 VDD VDD sg13_lv_pmos w=1u l=4u ng=1 m=1
XM5 net1 net3 VSS VSS sg13_lv_nmos w=2u l=2u ng=1 m=1
XM6 net3 net3 VSS VSS sg13_lv_nmos w=2u l=2u ng=1 m=1
I0 VDD net3 100n
.ends

.GLOBAL GND
.end
