** sch_path: /home/designer/shared/amaru/analog/tb/tb_rect_01.sch
**.subckt tb_rect_01
V1 VA VB dc 0 sin(0 500m 433Meg)
C1 VO1 VSS 100f m=1
V2 VSS GND 0
x1 VA VSS VO1 VB rect_01_10k
C2 VO2 VSS 100f m=1
x2 VA VO1 VO2 VB rect_01_10k
C3 VO3 VSS 100f m=1
x3 VA VO2 VO3 VB rect_01_10k
x4 VA VO3 VOUT VB rect_01_10k
C6 VOUT VSS 100f m=1
R1 net1 VSS 20k m=1
V3 VOUT net1 0
**** begin user architecture code


.param temp=27
.tran 0.1n 50u
.save VA VB VO1 VO2 VO3 VOUT I(V1) I(V3)
+ @n.x1.xm1.nsg13_lv_nmos[ids] @n.x1.xm2.nsg13_lv_nmos[ids]
+ @n.x1.xm3.nsg13_lv_pmos[ids] @n.x1.xm4.nsg13_lv_pmos[ids]
+ @n.x4.xm1.nsg13_lv_nmos[ids] @n.x4.xm2.nsg13_lv_nmos[ids]
+ @n.x4.xm3.nsg13_lv_pmos[ids] @n.x4.xm4.nsg13_lv_pmos[ids]

.control
  run
  let id1m1 = @n.x1.xm1.nsg13_lv_nmos[ids]
  let id1m2 = @n.x1.xm2.nsg13_lv_nmos[ids]
  let id1m3 = @n.x1.xm3.nsg13_lv_pmos[ids]
  let id1m4 = @n.x1.xm4.nsg13_lv_pmos[ids]
  let id4m1 = @n.x1.xm1.nsg13_lv_nmos[ids]
  let id4m2 = @n.x1.xm2.nsg13_lv_nmos[ids]
  let id4m3 = @n.x1.xm3.nsg13_lv_pmos[ids]
  let id4m4 = @n.x1.xm4.nsg13_lv_pmos[ids]
  write tb_rect_01.raw v(VA) v(VB) v(VO1) v(VO2) v(VO3) v(VOUT) I(V1) I(V3) id1m1 id1m2 id1m3 id1m4 id4m1 id4m2 id4m3 id4m4
.endc




.lib cornerMOSlv.lib mos_tt


**** end user architecture code
**.ends

* expanding   symbol:  rect_01_10k.sym # of pins=4
** sym_path: /home/designer/shared/amaru/analog/core/rect_01_10k.sym
** sch_path: /home/designer/shared/amaru/analog/core/rect_01_10k.sch
.subckt rect_01_10k VA VL VH VB
*.iopin VL
*.iopin VH
*.iopin VA
*.iopin VB
XM1 VL net1 net2 VL sg13_lv_nmos w=200u l=0.13u ng=40 m=1
XM3 VH net2 net1 VH sg13_lv_pmos w=400u l=0.13u ng=40 m=1
XM2 VL net2 net1 VL sg13_lv_nmos w=200u l=0.13u ng=40 m=1
XM4 VH net1 net2 VH sg13_lv_pmos w=400u l=0.13u ng=40 m=1
C1 VA net1 50p m=1
C2 net2 VB 50p m=1
.ends

.GLOBAL GND
.end
