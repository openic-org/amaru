** sch_path: /home/designer/shared/amaru/analog/core/inv_1x.sch
.subckt inv_1x VDD A Z VSS
*.PININFO VDD:B VSS:B A:B Z:B
M1 Z A VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M2 Z A VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
.ends
